module motion(
	input clk,
	input sense,
	output out
);


endmodule